
module Switches(din,dout);
    input [31:0] din;
	output [31:0] dout;
	
	//assign dout = din;
	assign dout = din;
endmodule